* /Users/marek/Documents/KiCad/debounced-clock/debounced-clock.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 2017 April 22, Saturday 21:38:17

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
R3  23 2 1K		
R7  18 1 220		
C5  22 1 0.1uF		
C4  21 1 0.01uF		
XU4  1 23 15 2 21 22 22 2 NE555		
R1  20 13 1K		
R2  20 2 1K		
C3  17 1 1uF		
C1  19 1 0.01uF		
P1  2 1 POWER		
XU1  1 17 12 2 19 17 20 2 NE555		
C2  2 1 0.01uF		
R4  2 22 1M		
C6  25 1 0.01uF		
XU5  1 9 4 24 25 1 ? 2 NE555		
P3  1 23 STEP		
P4  24 1 9 SWITCH		
P6  14 18 LED		
R5  9 2 1K		
R6  2 24 1K		
XU2  12 4 11 4 4 10 1 3 10 15 ? 16 16 2 7400		
XU3  11 3 6 6 ? 8 1 14 8 8 2 7400		
P5  16 HALT		
P7  2 1 POWER		
C7  2 1 0.01uF		
P2  13 17 POT		

.end
